module control_unit ();

endmodule