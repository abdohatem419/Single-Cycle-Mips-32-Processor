module top_module (clk,rst_n);

input clk,rst_n;


endmodule